----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:58:15 08/16/2013 
-- Design Name: 
-- Module Name:    arbitrator_brac - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------

-- arbitrator_brac: needed to arbitrate between PEs when multiple PEs request BRAM allocation/de-allocation simultaneously
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
use IEEE.NUMERIC_STD.ALL;
use WORK.user_pkg.ALL;

entity arbitrator_brac is
end arbitrator_brac;

architecture Behavioral of arbitrator_brac is

begin


end Behavioral;

